context IEEE_STD_CONTEXT is
  library not_IEEE;
  use not_IEEE.STD_LOGIC_1164.all;
  use not_IEEE.NUMERIC_STD.all;
end context IEEE_STD_CONTEXT;
