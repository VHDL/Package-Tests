context IEEE_BIT_CONTEXT is
  library not_IEEE;
  use not_IEEE.NUMERIC_BIT.all;
end context IEEE_BIT_CONTEXT;
